module spi_tb (
);
    
endmodule