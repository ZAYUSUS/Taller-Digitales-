
module Spi (
    ports
);


endmodule