
module TB;
ALU alu0();
endmodule